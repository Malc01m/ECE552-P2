module MEM_WB_buf();
endmodule