module EX_MEM_buf();
endmodule