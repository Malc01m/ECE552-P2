module hazardUnit();
endmodule